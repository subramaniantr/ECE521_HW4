vin 1 0 5
r1 1 2 2000
d1 2 3 dmod 1
r2 3 0 3000
