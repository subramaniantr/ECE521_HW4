vcc 1 0 5
rc1 1 2 1000
q1 2 3 0 npn
r12 3 4 500
rc2 1 5 500
q2 5 4 6 npn
re2 6 0 500
vb 3 0 0.78
